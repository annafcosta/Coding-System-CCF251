module moduleConv (
    By1, By2, By3, By4,
    s0, s1, s2, s3
    ready, reset
);
input wire By1;
input wire By2;
input wire By3;
input wire By4;



output reg s0;
output reg s1;
output reg s2;
output reg s3;

    
endmodule