/*module lot_tb;
	reg clk_tb, reset_tb, fim_tb, fim_jogo_tb, insere_tb;
	reg [0:3] num_tb;
	wire [0:1] premio_tb;
	wire [0:4] p1_tb, p2_tb;

	Lot TB (.clk(clk_tb), .reset(reset_tb), .fim(fim_tb), .fim_jogo(fim_jogo_tb), .insere(insere_tb),
				.num(num_tb), .premio(premio_tb), .p1(p1_tb), .p2(p2_tb));
				
	initial begin
		
		$dumpfile("teste_gtx.vcd");
		$dumpvars;
	
	
	
		clk_tb = 0;
		reset_tb = 1;
		fim_tb = 0;
		fim_jogo_tb = 0;
		insere_tb = 0;
		
		
		
		
		
		
		
		
		
		
		
		
		
		
	end
	


endmodule */
