module HelloWorld;

  initial begin
    $display("Hello, World!");
    $finish;
  end

endmodule
